module conv (input W, X, Y, Z, output outa,outb,outc,outd,oute,outf,outg );

a a1(W, X, Y, Z,outa);
b b1(W, X, Y, Z,outb);
c c1(W, X, Y, Z,outc);
d d1(W, X, Y, Z,outd);
e e1(W, X, Y, Z,oute);
f f1(W, X, Y, Z,outf);
g g1(W, X, Y, Z,outg);

endmodule


